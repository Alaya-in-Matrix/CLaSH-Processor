// Automatically generated Verilog-2001
module System_testInput_11(topLet_o);
  output [16:0] topLet_o;
  assign topLet_o = {1'b1
                    ,16'sd2};
endmodule
